library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.epu_pack.all;

entity prom is
	port(
		I_Addr	: in std_logic_vector(3 downto 0);
		O_M		: out std_logic_vector(0 to 31)
	);
end prom;

architecture prom_behav of prom is
	type rom_array is array (NATURAL range <>) of std_logic_vector(0 to 31);

	constant rom : rom_array := (
		"01111111111011111111101000000010",
		"01000000000010000000101000000010",
		"01000000000010000000101000000010",
		"01000000000010000000101000000010",
		"01000000000010000000101000000010",
		"01000000000010000000101000000010",
		"01000000000011111111101000000010",
		"01111111111010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01000000000010000000001000000010",
		"01111111111010000000001111111110"
	);
begin
	process(I_Addr)
	begin
		O_M <= rom(to_integer(unsigned(I_Addr)));
	end process;
end prom_behav;
